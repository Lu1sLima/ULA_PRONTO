library IEEE;
use IEEE.Std_Logic_1164.all;
package p_ula is
type op_alu is
( uAND, uOR, uXNOR, uSLL, uSRL, uADD, uSUB, uSUB2, uOP1, uNEG);
end p_ula;
